// ======================================================
//                      VI SEnC 2022
// ======================================================

module MercurioIV_nios_top(

    //////// CLOCK //////////
    CLOCK_50MHz,

    //////// LED //////////
    LEDM_C,
    LEDM_R,

    //////// KEY //////////
    KEY,

    //////// SW //////////
    SW
);

//=======================================================
//  PARAMETER declarations
//=======================================================


//=======================================================
//  PORT declarations
//=======================================================

//////////// CLOCK //////////
input                    CLOCK_50MHz;

//////////// LED //////////
output         [4:0]     LEDM_C;
output         [7:0]     LEDM_R;

//////////// KEY //////////
input          [11:0]     KEY;

//////////// SW //////////
input          [3:0]     SW;

/////////////////////////////////////////////////////////
//=======================================================
// REG/WIRE declarations
//=======================================================


//=======================================================
// Structural coding
//=======================================================

assign	LEDM_C        =    5'bz;
assign	LEDM_R        =    8'bz;

endmodule
