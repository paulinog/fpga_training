// ======================================================
//                      VI SEnC 2022
// ======================================================

module MercurioIV_fsm_top(

    //////// CLOCK //////////
    CLOCK_50MHz,

    //////// LED //////////
    LEDM_C,
    LEDM_R,

    //////// KEY //////////
    KEY
);

//=======================================================
//  PARAMETER declarations
//=======================================================


//=======================================================
//  PORT declarations
//=======================================================

//////////// CLOCK //////////
input                    CLOCK_50MHz;

//////////// LED //////////
output         [4:0]     LEDM_C;
output         [7:0]     LEDM_R;

//////////// KEY //////////
input          [11:0]     KEY;

/////////////////////////////////////////////////////////
//=======================================================
// REG/WIRE declarations
//=======================================================


//=======================================================
// Structural coding
//=======================================================

assign	LEDM_C        =    5'bz;
assign	LEDM_R        =    8'bz;

// mealy_mac u2
// (
// 	.clk(CLOCK_50), 
// 	.data_in(KEY[1]), 
// 	.reset(KEY[0]),
// 	.data_out(LEDM_R[1:0])
// );

endmodule
